`timescale 1ns/1ns
`include "question1b.v"

module question1b_tb();
  reg a,b,c,d;
  wire f;

  question1b q1b(a,b,c,d,f);
  initial 
    begin 
      $dumpfile("question1b_tb.vcd");
      $dumpvars(0,question1b_tb);

      a=1'b0; b=1'b0; c=1'b0; d=1'b0;
      #20
      a=1'b0; b=1'b0; c=1'b0; d=1'b1;
      #20
      a=1'b0; b=1'b0; c=1'b1; d=1'b0;
      #20
      a=1'b0; b=1'b0; c=1'b1; d=1'b1;
      #20
      a=1'b0; b=1'b1; c=1'b0; d=1'b0;
      #20
      a=1'b0; b=1'b1; c=1'b0; d=1'b1;
      #20
      a=1'b0; b=1'b1; c=1'b1; d=1'b0;
      #20
      a=1'b0; b=1'b1; c=1'b1; d=1'b1;
      #20
      a=1'b1; b=1'b0; c=1'b0; d=1'b0;
      #20
      a=1'b1; b=1'b0; c=1'b0; d=1'b1;
      #20
      a=1'b1; b=1'b0; c=1'b1; d=1'b0;
      #20
      a=1'b1; b=1'b0; c=1'b1; d=1'b1;
      #20
      a=1'b1; b=1'b1; c=1'b0; d=1'b0;
      #20
      a=1'b1; b=1'b1; c=1'b0; d=1'b1;
      #20
      a=1'b1; b=1'b1; c=1'b1; d=1'b0;
      #20
      a=1'b1; b=1'b1; c=1'b1; d=1'b1;
      #20

      $display("Test Complete");
    end
endmodule